-- Libraries
library ieee;
use ieee.std_logic_1164.all;

-- Chapter 4 - Example 4