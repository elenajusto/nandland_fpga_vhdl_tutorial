-- File: Top Level

-- ***** Project Entities *****

-- Definition: 1 Hz Counter

-- Definition: 10 Hz Counter

-- Definition: 50 Hz Counter

-- Definition: 100 Hz Counter

-- Definition: Switch 1

-- Definition: Switch 2

-- Definition: Enable

-- Definition: Multiplixer

-- Definition: AND Gate

-- ***** Project Interaction *****
-- 1 Hz clock signal entering 1 Hz counter
-- 10 Hz clock signal entering 10 Hz counter
-- 50 Hz clock signal entering 50 Hz counter
-- 100 Hz clock signal entering 100 Hz counter