-- Libraries
library ieee;
use ieee.std_logic_1164.all;

-- Chapter 4 - Example 7
-- Write the VHDL code that implements the following  circuit. 
-- The circuit contains an input bundle of four signals and
-- an output bundle of three signals. 
-- The input bundle, D IN, represents a 4bit binary number. 
-- The output bundle, SZ OUT, is used to indicate the magnitude 
-- of the 4-bit binary input number. 

-- The relationship between  the input and output is shown in 
-- the table below. 

-- Use a selected signal  assignment statement in the solution.
